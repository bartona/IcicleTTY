----------------------------------------------------------------------
-- Created by Actel SmartDesign Tue Oct 01 22:52:07 2013
-- Parameters for COREUART
----------------------------------------------------------------------


package coreparameters is
    constant BAUD_VAL_FRCTN_EN : integer := 0;
    constant FAMILY : integer := 20;
    constant HDL_license : string( 1 to 1 ) := "O";
    constant RX_FIFO : integer := 0;
    constant RX_LEGACY_MODE : integer := 0;
    constant testbench : string( 1 to 4 ) := "User";
    constant TX_FIFO : integer := 0;
    constant USE_SOFT_FIFO : integer := 0;
end coreparameters;
